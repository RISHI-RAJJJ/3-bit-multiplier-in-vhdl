library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_arith.all;
entity multt is
port(b0,b1,b2,a0,a1,a2 :in std_logic;
     p0,p1,p2,p3,p4,p5,p6,c1,s1,c2,c3,c4,c5,c6,c7,s2,s3 :out std_logic);
end multt ;

architecture multt of multt is
begin
p0 <= (b0 and a0) ;
p1 <= ((b0 and a1) xor (b1 and a0) xor '0');
c1 <= (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'));
s1 <= ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')));
c3 <= (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))));
p2 <= ('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))) xor (b2 and a0));
c2 <= (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)));
s2 <= ('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))));
c4 <= (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))));
p3 <= (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) xor (b1 and a2) xor (b2 and a1));
c5 <= ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) and (b1 and a2)) or ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) xor (b1 and a2)) and (b2 and a1)));
s3 <= ('0' xor (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))))) xor ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) and (b1 and a2)) or ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) xor (b1 and a2)) and (b2 and a1))));
c6 <= (('0' and (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))))) or (('0' xor (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))))) and ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) and (b1 and a2)) or ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) xor (b1 and a2)) and (b2 and a1)))));
p4 <= ('0' xor (b2 and a2) xor ('0' xor (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))))) xor ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) and (b1 and a2)) or ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) xor (b1 and a2)) and (b2 and a1)))));
c7 <= (('0' and (b2 and a2)) or (('0' xor (b2 and a2)) and ('0' xor (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))))) xor ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) and (b1 and a2)) or ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) xor (b1 and a2)) and (b2 and a1))))));
p5 <= ('0' xor (('0' and (b2 and a2)) or (('0' xor (b2 and a2)) and ('0' xor (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))))) xor ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) and (b1 and a2)) or ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) xor (b1 and a2)) and (b2 and a1)))))) xor (('0' and (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))))) or (('0' xor (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))))) and ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) and (b1 and a2)) or ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) xor (b1 and a2)) and (b2 and a1))))));
p6 <= (('0' and (('0' and (b2 and a2)) or (('0' xor (b2 and a2)) and ('0' xor (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))))) xor ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) and (b1 and a2)) or ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) xor (b1 and a2)) and (b2 and a1))))))) or (('0' xor (('0' and (b2 and a2)) or (('0' xor (b2 and a2)) and ('0' xor (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))))) xor ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) and (b1 and a2)) or ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) xor (b1 and a2)) and (b2 and a1))))))) and (('0' and (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))))) or (('0' xor (('0' and (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) or (('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0)))) and (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))))) and ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) and (b1 and a2)) or ((('0' xor (('0' and ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) or (('0' xor ((b1 and a1) xor (b0 and a2) xor (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0')))) and (b2 and a0))) xor (((b1 and a1) and (b0 and a2)) or (((b1 and a1) xor (b0 and a2)) and (((b0 and a1) and (b1 and a0)) or (((b0 and a1) xor (b1 and a0)) and '0'))))) xor (b1 and a2)) and (b2 and a1)))))));
end multt ;